/*`define MINUSONE_ 110
`define MINUSTWO_ 101
`define ZERO_ 	  000
`define ONE_	  001
`define TWO_	  010
 */
module quotient_selection
		#(parameter ND=4,
			    NP=7 //3bits after decimal and 4 before decimal 0000.000
		 )		
		(input [ND-1:0]d,  //the divisor as x cordinate
		       [NP-1:0]rpj, //the shifted partial remainder as y cordinate			
		 output reg[2:0] q_jplus1 //q[j+1] in rbsd form		
		);
	
reg [47:0] temp_row;

always @(rpj)begin
case(rpj)
		
	7'b0101011: temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_010;

	7'b0101010: temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_010_010;

	7'b0101001: temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_010_010;
	
	7'b0101000:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_010_010_010;

	7'b0100111:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_010_010_010_010;

	7'b0100110:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_010_010_010_010_010;

	7'b0100101:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_010_010_010_010_010;

	7'b0100100:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_010_010_010_010_010_010;

	7'b0100011:temp_row = 48'b000_000_000_000_000_000_000_000_000_010_010_010_010_010_010_010;

	7'b0100010:temp_row = 48'b000_000_000_000_000_000_000_000_000_010_010_010_010_010_010_010;

	7'b0100001:temp_row = 48'b000_000_000_000_000_000_000_000_010_010_010_010_010_010_010_010;

	7'b0100000:temp_row = 48'b000_000_000_000_000_000_000_010_010_010_010_010_010_010_010_010;

	7'b0011111:temp_row = 48'b000_000_000_000_000_000_010_010_010_010_010_010_010_010_010_010;

	7'b0011110:temp_row = 48'b000_000_000_000_000_010_010_010_010_010_010_010_010_010_010_010;

	7'b0011101:temp_row = 48'b000_000_000_000_000_010_010_010_010_010_010_010_010_010_010_010;

	7'b0011100:temp_row = 48'b000_000_000_000_010_010_010_010_010_010_010_010_010_010_010_010;

	7'b0011011:temp_row = 48'b000_000_000_010_010_010_010_010_010_010_010_010_010_010_010_010;

	7'b0011010:temp_row = 48'b000_000_010_010_010_010_010_010_010_010_010_010_010_010_010_010;

	7'b0011001:temp_row = 48'b000_000_010_010_010_010_010_010_010_010_010_010_010_010_010_010;

	7'b0011000:temp_row = 48'b000_010_010__010_010_010_010_010_010_010_010_010_010_010_010_010;
	
	7'b0010111:temp_row = 48'b010_010_010_010_010_010_010_010_010_010_010_010_010_010_010_010;
	
	7'b0010110:temp_row = 48'b010_010_010_010_010_010_010_010_010_010_010_010_010_010_001_001;
	
	7'b0010101:temp_row = 48'b010_010_010_010_010_010_010_010_010_010_010_010_010_010_001_001;
	
	7'b0010100:temp_row = 48'b010_010_010_010_010_010_010_010_010_010_010_001_001_001_001_001;
	
	7'b0010011:temp_row = 48'b010_010_010_010_010_010_010_010_010_010_010_001_001_001_001_001;
	
	7'b0010010:temp_row = 48'b010_010_010_010_010_010_010_010_001_001_001_001_001_001_001_001;
	
	7'b0010001:temp_row = 48'b010_010_010_010_010_010_010_010_001_001_001_001_001_001_001_001;
	
	7'b0010000:temp_row = 48'b010_010_010_010_010_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001111:temp_row = 48'b010_010_010_010_010_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001110:temp_row = 48'b010_010_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001101:temp_row = 48'b010_010_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001100:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001011:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001010:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001001:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0001000:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0000111:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_001_001;
	
	7'b0000110:temp_row = 48'b001_001_001_001_001_001_001_001_001_001_001_001_001_001_000_000;
	
	7'b0000101:temp_row = 48'b001_001_001_001_001_001_001_001_000_000_000_000_000_000_000_000;
	
	7'b0000100:temp_row = 48'b001_001_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b0000011:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b0000010:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b0000001:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b0000000:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b1111111:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b1111110:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b1111101:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b1111100:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b1111011:temp_row = 48'b110_110_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
	
	7'b1111010:temp_row = 48'b110_110_110_110_110_110_110_110_000_000_000_000_000_000_000_000;
	
	7'b1111001:temp_row = 48'b110_110_110_110_110_110_110_110_110_110_110_110_110_110_000_000;
			
	7'b1111000:temp_row = 48'b110_110_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
			
	7'b1110111:temp_row = 48'b110_110_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
		
	7'b1110110:temp_row = 48'b110_110_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
		
	7'b1110101:temp_row = 48'b110_110_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
	
	7'b1110100:temp_row = 48'b110_110_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
	
	7'b1110011:temp_row = 48'b101_101_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
	
	7'b1110010:temp_row = 48'b101_101_110_110_110_110_110_110_110_110_110_110_110_110_110_110;
	
	7'b1110001:temp_row = 48'b101_101_101_101_010_110_110_110_110_110_110_110_110_110_110_110;
	
	7'b1110000:temp_row = 48'b101_101_101_101_101_110_110_110_110_110_110_110_110_110_110_110;
	
	7'b1101111:temp_row = 48'b101_101_101_101_101_101_101_101_110_110_110_110_110_110_110_110;
	
	7'b1101110:temp_row = 48'b101_101_101_101_101_101_101_101_110_110_110_110_110_110_110_110;
	
	7'b1101101:temp_row = 48'b101_101_101_101_101_101_101_101_101_101_101_110_110_110_110_110;
	
	7'b1101100:temp_row = 48'b101_101_101_101_101_101_101_101_101_101_101_110_110_110_110_110;
	
	7'b1101011:temp_row = 48'b101_101_101_101_101_101_101_101_101_101_101_101_101_101_110_110;
	
	7'b1101010:temp_row = 48'b101_101_101_101_101_101_101_101_101_101_101_101_101_101_110_110;
	
	7'b1101001:temp_row = 48'b000_101_101_101_101_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1101000:temp_row = 48'b000_000_101_101_101_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100111:temp_row = 48'b000_000_101_101_101_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100110:temp_row = 48'b000_000_000_101_101_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100101:temp_row = 48'b000_000_000_000_101_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100100:temp_row = 48'b000_000_000_000_000_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100011:temp_row = 48'b000_000_000_000_000_101_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100010:temp_row = 48'b000_000_000_000_000_000_101_101_101_101_101_101_101_101_101_101;
	
	7'b1100001:temp_row = 48'b000_000_000_000_000_000_000_000_000_101_101_101_101_101_101_101;
	
	7'b1100000:temp_row = 48'b000_000_000_000_000_000_000_000_101_101_101_101_101_101_101_101;
	
	7'b1011111:temp_row = 48'b000_000_000_000_000_000_000_000_101_101_101_101_101_101_101_101;
	
	7'b1011110:temp_row = 48'b000_000_000_000_000_000_000_000_000_101_101_101_101_101_101_101;
	
	7'b1011101:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_101_101_101_101_101_101;
	
	7'b1011100:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_101_101_101_101_101;
	
	7'b1011011:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_101_101_101_101_101;
	
	7'b1011010:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_101_101_101_101;
	
	7'b1011001:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_101_101_101;
	
	7'b1011000:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_101_101;
	
	7'b1010111:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_101_101;
	
	7'b1010110:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_101;
	
	7'b1010101:temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_101;	
	
	default : temp_row = 48'b000_000_000_000_000_000_000_000_000_000_000_000_000_000_000_000;
		
	endcase
end

always @(d, temp_row) begin
	case (d) 
		4'b1111 : q_jplus1 = temp_row[2:0];
		
		4'b1110 : q_jplus1 = temp_row[5:3];
		
		4'b1101 : q_jplus1 = temp_row[8:6];
	
		4'b1100 : q_jplus1 = temp_row[11:9];
		
		4'b1011 : q_jplus1 = temp_row[14:12];
		
		4'b1010 : q_jplus1 = temp_row[17:15];
		
		4'b1001 : q_jplus1 = temp_row[20:18];
		
		4'b1000 : q_jplus1 = temp_row[23:21];
		
		4'b0111 : q_jplus1 = temp_row[26:24];
		
		4'b0110 : q_jplus1 = temp_row[39:27];
		
		4'b0101 : q_jplus1 = temp_row[32:30];
		
		4'b0100 : q_jplus1 = temp_row[35:33];
	
		4'b0011 : q_jplus1 = temp_row[38:36];
		
		4'b0010 : q_jplus1 = temp_row[41:39];
		
		4'b0001 : q_jplus1 = temp_row[44:42];
		
		4'b0000 : q_jplus1 = temp_row[47:45];
		
	endcase
end

endmodule
/*
module top;
reg [3:0]d;
reg [6:0]rpj;
wire [2:0]q_jplus1;

	quotient_selection qs1(d,rpj,q_jplus1);

initial begin
	d = 4'b1100;
	rpj = 7'b1111_100;
end

initial begin
	$monitor("d = %b, rpj = %b, \n temp_row = %b, q_jplus1 = %b",d,rpj,qs1.temp_row,q_jplus1);
end
endmodule
*/